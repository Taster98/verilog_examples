module not_m(output z, input x);
    //qui faccio tutti gli assegnamenti
    assign
        z = ~x;
endmodule